magic
tech sky130A
timestamp 1714035034
<< nwell >>
rect -150 -150 150 300
<< nmos >>
rect -10 -300 5 -200
<< pmos >>
rect -10 -100 5 105
<< ndiff >>
rect -55 -210 -10 -200
rect -55 -290 -45 -210
rect -25 -290 -10 -210
rect -55 -300 -10 -290
rect 5 -210 50 -200
rect 5 -290 20 -210
rect 40 -290 50 -210
rect 5 -300 50 -290
<< pdiff >>
rect -60 95 -10 105
rect -60 -95 -50 95
rect -25 -95 -10 95
rect -60 -100 -10 -95
rect 5 95 55 105
rect 5 -95 20 95
rect 45 -95 55 95
rect 5 -100 55 -95
<< ndiffc >>
rect -45 -290 -25 -210
rect 20 -290 40 -210
<< pdiffc >>
rect -50 -95 -25 95
rect 20 -95 45 95
<< psubdiff >>
rect -60 -355 55 -340
rect -60 -380 -45 -355
rect 40 -380 55 -355
rect -60 -395 55 -380
<< nsubdiff >>
rect -95 250 90 265
rect -95 220 -80 250
rect 75 220 90 250
rect -95 205 90 220
<< psubdiffcont >>
rect -45 -380 40 -355
<< nsubdiffcont >>
rect -80 220 75 250
<< poly >>
rect -10 105 5 165
rect -10 -200 5 -100
rect -10 -330 5 -300
<< locali >>
rect -95 250 90 265
rect -95 220 -80 250
rect 75 220 90 250
rect -95 205 90 220
rect -60 95 -15 105
rect -60 -95 -50 95
rect -25 -95 -15 95
rect -60 -100 -15 -95
rect 10 95 55 105
rect 10 -95 20 95
rect 45 -95 55 95
rect 10 -100 55 -95
rect -55 -210 -15 -200
rect -55 -290 -45 -210
rect -25 -290 -15 -210
rect -55 -300 -15 -290
rect 10 -210 50 -200
rect 10 -290 20 -210
rect 40 -290 50 -210
rect 10 -300 50 -290
rect -55 -355 50 -345
rect -55 -380 -45 -355
rect 40 -380 50 -355
rect -55 -390 50 -380
<< end >>
