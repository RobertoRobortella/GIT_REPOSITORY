magic
tech sky130A
timestamp 1714038282
<< nwell >>
rect -150 -150 150 300
<< nmos >>
rect -10 -300 5 -200
<< pmos >>
rect -10 -100 5 105
<< ndiff >>
rect -55 -210 -10 -200
rect -55 -290 -45 -210
rect -25 -290 -10 -210
rect -55 -300 -10 -290
rect 5 -210 50 -200
rect 5 -290 20 -210
rect 40 -290 50 -210
rect 5 -300 50 -290
<< pdiff >>
rect -60 95 -10 105
rect -60 -95 -50 95
rect -25 -95 -10 95
rect -60 -100 -10 -95
rect 5 95 55 105
rect 5 -95 20 95
rect 45 -95 55 95
rect 5 -100 55 -95
<< ndiffc >>
rect -45 -290 -25 -210
rect 20 -290 40 -210
<< pdiffc >>
rect -50 -95 -25 95
rect 20 -95 45 95
<< psubdiff >>
rect -95 -355 100 -340
rect -95 -375 -80 -355
rect 85 -375 100 -355
rect -95 -390 100 -375
<< nsubdiff >>
rect -95 250 90 265
rect -95 220 -80 250
rect 75 220 90 250
rect -95 205 90 220
<< psubdiffcont >>
rect -80 -375 85 -355
<< nsubdiffcont >>
rect -80 220 75 250
<< poly >>
rect -10 105 5 165
rect -10 -140 5 -100
rect -85 -150 5 -140
rect -85 -170 -75 -150
rect -45 -170 5 -150
rect -85 -180 5 -170
rect -10 -200 5 -180
rect -10 -330 5 -300
<< polycont >>
rect -75 -170 -45 -150
<< locali >>
rect -95 255 90 265
rect -95 250 -30 255
rect 15 250 90 255
rect -95 220 -80 250
rect 75 220 90 250
rect -95 215 -30 220
rect 15 215 90 220
rect -95 205 90 215
rect -60 95 -15 205
rect -60 -95 -50 95
rect -25 -95 -15 95
rect -60 -100 -15 -95
rect 10 95 55 105
rect 10 -95 20 95
rect 45 -95 55 95
rect 10 -140 55 -95
rect -85 -150 -25 -140
rect -85 -170 -75 -150
rect -45 -170 -25 -150
rect -85 -180 -25 -170
rect 10 -150 125 -140
rect 10 -170 90 -150
rect 115 -170 125 -150
rect 10 -180 125 -170
rect -55 -210 -15 -200
rect -55 -290 -45 -210
rect -25 -290 -15 -210
rect -55 -340 -15 -290
rect 10 -210 55 -180
rect 10 -290 20 -210
rect 40 -275 55 -210
rect 40 -290 50 -275
rect 10 -300 50 -290
rect -95 -350 100 -340
rect -95 -355 -55 -350
rect 45 -355 100 -350
rect -95 -375 -80 -355
rect 85 -375 100 -355
rect -95 -385 -55 -375
rect 45 -385 100 -375
rect -95 -390 100 -385
rect -55 -395 -15 -390
<< viali >>
rect -30 250 15 255
rect -30 220 15 250
rect -30 215 15 220
rect -75 -170 -45 -150
rect 90 -170 115 -150
rect -55 -355 45 -350
rect -55 -375 45 -355
rect -55 -385 45 -375
<< metal1 >>
rect -325 255 335 265
rect -325 215 -30 255
rect 15 215 335 255
rect -325 205 335 215
rect -355 -150 -25 -140
rect -355 -170 -75 -150
rect -45 -170 -25 -150
rect -355 -180 -25 -170
rect 10 -150 340 -140
rect 10 -170 90 -150
rect 115 -170 340 -150
rect 10 -190 340 -170
rect -320 -350 340 -335
rect -320 -385 -55 -350
rect 45 -385 340 -350
rect -320 -395 340 -385
<< labels >>
rlabel metal1 255 230 255 230 1 vdd
rlabel metal1 230 -365 230 -365 1 vss
rlabel metal1 280 -170 305 -160 1 out
rlabel metal1 -335 -165 -310 -155 1 in
<< end >>
